//MDR