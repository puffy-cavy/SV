//IR