//MAR
